module multiplier (input a,
	input b,
	output p);
	assign p=a*b;
endmodule
